----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Fu Zuoyou.
-- 
-- Create Date:    17:12:10 11/26/2013 
-- Design Name: 
-- Module Name:    VGA_play - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity VGA_play is
	Port(
		CLK_0: in std_logic;
		reset: in std_logic;
		R: out std_logic_vector(2 downto 0) := "000";
		G: out std_logic_vector(2 downto 0) := "000";
		B: out std_logic_vector(2 downto 0) := "000";
		Hs: out std_logic := '0';
		Vs: out std_logic := '0';
		hclk: in std_logic
	);
end VGA_play;

architecture Behavioral of VGA_play is
	signal clk: std_logic;
	signal vector_x : std_logic_vector(9 downto 0);		--X 640
	signal vector_y : std_logic_vector(8 downto 0);		--Y 480
	signal r0 : std_logic_vector(2 downto 0);
	signal g0 : std_logic_vector(2 downto 0);
	signal b0 : std_logic_vector(2 downto 0);
	signal hs1 : std_logic;
	signal vs1 : std_logic;

	signal char: std_logic_vector(7 downto 0) := "00000000";
	signal pr: std_logic_vector(7 downto 0);
	signal tmpp: std_logic_vector(11 downto 0);
	
	component char_mem
	  PORT (
		clka : IN STD_LOGIC;
		addra : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		douta : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	  );
	end component;
	signal tmp2: std_logic_vector (3 downto 0);
begin

	ram: char_mem port map(clka => clk, addra => tmpp, douta => pr);
	
	tmpp <=  char(7 downto 0) & vector_y(8 downto 5);
	tmp2 <= vector_x(3 downto 0);

process(hclk)
begin
	if hclk'event and hclk = '1' then
		char <= char + 1;
	end if;
end process;

-- 50 MHz -> 25 MHz
process(CLK_0)
begin
	if(CLK_0'event and CLK_0 = '1') then
		clk <= not clk;
	end if;
end process;

process(clk, reset)	-- ������������ (800)
begin
	if reset = '0' then
		vector_x <= (others => '0');
	elsif clk'event and clk = '1' then
		if vector_x = 799 then
			vector_x <= (others => '0');
		else
			vector_x <= vector_x + 1;
		end if;
	end if;
end process;

process(clk, reset)	-- ���������� (525)
begin
	if reset = '0' then
		vector_y <= (others => '0');
	elsif clk'event and clk = '1' then
		if vector_x = 799 then
			if vector_y = 524 then
				vector_y <= (others => '0');
			else
				vector_y <= vector_y + 1;
			end if;
		end if;
	end if;
end process;

process(clk, reset) -- ��ͬ���źţ�640+��������16��+96��+48�գ�
begin
	if reset='0' then
		hs1 <= '1';
	elsif clk'event and clk='1' then
		if vector_x >= 656 and vector_x < 752 then
			hs1 <= '0';
		else
			hs1 <= '1';
		end if;
	end if;
end process;

process(clk, reset) -- ��ͬ���źţ�480+��������10��+2��+33�գ�
begin
	if reset = '0' then
		vs1 <= '1';
	elsif clk'event and clk = '1' then
		if vector_y >= 490 and vector_y < 492 then
			vs1 <= '0';
		else
			vs1 <= '1';
		end if;
	end if;
end process;

process(clk, reset)
begin
	if reset = '0' then
		hs <= '0';
		vs <= '0';
	elsif clk'event and clk = '1' then
		hs <= hs1;
		vs <= vs1;
	end if;
end process;

process(reset, clk, vector_x, vector_y) -- X, Y �������
begin
	if reset = '0' then
		r0 <= "000";
		g0 <= "000";
		b0 <= "000";
	elsif clk'event and clk = '1' then
		if vector_x > 639 or vector_y > 479 then
			r0 <= "000";
			g0 <= "000";
			b0 <= "000";
		else		
			-- play around
			if tmp2 >= 0 and tmp2 < 2 then			
				if pr(0) = '1' then
					r0 <= "111";g0 <= "000";b0 <= "000";
				else
					r0 <= "000";g0 <= "000";b0 <= "000";
				end if;
			elsif tmp2 >= 2 and tmp2 < 4 then			
				if pr(1) = '1'  then
					r0 <= "111";g0 <= "000";b0 <= "000";
				else
					r0 <= "000";g0 <= "000";b0 <= "000";
				end if;
			elsif tmp2 >= 4 and tmp2 < 6 then			
				if pr(2)  = '1' then
					r0 <= "111";g0 <= "000";b0 <= "000";
				else
					r0 <= "000";g0 <= "000";b0 <= "000";
				end if;
			elsif tmp2 >= 6 and tmp2 < 8 then			
				if pr(3)  = '1' then
					r0 <= "111";g0 <= "000";b0 <= "000";
				else
					r0 <= "000";g0 <= "000";b0 <= "000";
				end if;
			elsif tmp2 >= 8 and tmp2 < 10 then			
				if pr(4)  = '1' then
					r0 <= "111";g0 <= "000";b0 <= "000";
				else
					r0 <= "000";g0 <= "000";b0 <= "000";
				end if;
			elsif tmp2 >= 10 and tmp2 < 12 then			
				if pr(5)  = '1' then
					r0 <= "111";g0 <= "000";b0 <= "000";
				else
					r0 <= "000";g0 <= "000";b0 <= "000";
				end if;
			elsif tmp2 >= 12 and tmp2 < 14 then			
				if pr(6)  = '1' then
					r0 <= "111";g0 <= "000";b0 <= "000";
				else
					r0 <= "000";g0 <= "000";b0 <= "000";
				end if;
			elsif tmp2 >= 14 and tmp2 < 16 then			
				if pr(7)  = '1' then
					r0 <= "111";g0 <= "000";b0 <= "000";
				else
					r0 <= "000";g0 <= "000";b0 <= "000";
				end if;
			end if;
		end if;
	end if;
end process;

process(hs1, vs1, r0, g0, b0) -- ��͵�ɫ�����
begin
	if hs1 = '1' and vs1 = '1' then
		R <= r0;
		G <= g0;
		B <= b0;
	else
		R <= (others => '0');
		G <= (others => '0');
		B <= (others => '0');
	end if;
end process;

end Behavioral;

